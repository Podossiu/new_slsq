b0VIM 8.2      t�{c�k�� ilena7440                               eslab10                                 ~ilena7440/new/SLSQ_FINAL/quan/quantizer/lsq.py                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              utf-8 3210    #"! U                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 tp           j                            J       k                     ]       �                     c                                  u                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     ad  p   4     j       �  �  �  �  �  �  �  u  k  T  *  )  (      �  �  �  �  O  N  ;  )    �  �  �  �  q  P  5  ,      �  �  �  �  �  �  d  R  <  (  #    �  �  �  �  d    �
  �
  �
  �
  �
  k
  B
  A
  
  �	  �	  �	  |	  S	  '	  	  �  1  0  �  �  �  �  �  �  �  �  u  N  "  �  �  �  �  X  1  ,    �  �  4    �  �  �  �  �  �  2  �  �  �  V  4  3                                                                                                                          if not self.hard_pruning:         #score = x_reshape.abs().mean(dim = 1,keepdim = True)         score = x_reshape.abs().mean(dim = 1,keepdim = True) - p         #p = grad_scale(p, p_grad_scale)         #score = score / (score.max().detach() * 2)         x_reshape = x.reshape(co // self.block_size, self.block_size, ci, kh, kw)                  co, ci, kh, kw = x.shape      def soft_pruner(self, x, p):          return hard_mask.sum(), hard_mask.numel()         hard_mask = (score > 0).float().detach()         score = (x_reshape.abs().mean(dim = 1, keepdim = True) - self.p).detach()         x_reshape = x.reshape(co // self.block_size, self.block_size, ci, kh, kw).detach()         co, ci, kh, kw = x.shape     def calculate_block_sparsity(self,x):              self.temperature = temperature         self.hard_pruning = hard_pruning         self.block_size = block_size         self.soft_mask = None         self.weight_quantizer = weight_quant.apply         self.c = t.nn.Parameter(t.ones(1))         self.p= t.nn.Parameter(t.zeros([]))         self.per_channel = per_channel         self.thd_pos = 2 ** (bit - 1) - 1         self.thd_neg = -2 ** (bit - 1) + 1                  super().__init__(bit)     def __init__(self, bit, per_channel=False, symmetric = False, all_positive = False, hard_pruning = False, block_size = 4, temperature = 1e-3): class SLsqQuan(Quantizer):          return grad_input, grad_c, grad_p, None         #grad_input = ((1. - s_mask) + s_mask * thd * v_t * ste_constant) * grad_output.clone()          #grad_c = ((grad_c - s_mask * ste_constant * v_t * sign) * grad_output.clone()).sum().reshape(c.shape)         #grad_p = ((grad_p + s_mask * ste_constant * v_t * (-thd + 0.5) * sign) * grad_output.clone()).sum().reshape(p.shape)                  #ste_constant = 2 * s / (2 * p + s)         grad_input = grad_output.clone()         grad_p = (grad_p * grad_output.clone()).sum()         grad_c = (grad_c * grad_output.clone()).sum()                  grad_p = grad_p - sign * c_mask         grad_c = grad_c + sign * c_mask          grad_p = -grad_c - sign * i_mask         grad_c = (v_q / thd - v_t * sign) * i_mask                  v_t = (input.abs() - p) / distance                  sign = input.sign()         s_mask = (v_q == 0.).float()         i_mask =(input.abs() <= c).float() * (input.abs() >= p).float()         c_mask =(input.abs() > c).float()         thd = ctx.thd         s = ctx.s         input, v_q, c, p, distance = ctx.saved_tensors     def backward(ctx, grad_output):     @staticmethod              return v_dq         ctx.thd = thd         ctx.s = s         ctx.save_for_backward(input, v_q, c, p, distance)                  v_dq = v_q * s          v_q = t.round(v_c)          v_c = t.clamp(v_g, 0, thd) * sign            v_g = (input.abs() - p) / s                  s = distance / thd         distance = c - p + 1e-12         sign = input.sign()     def forward(ctx, input, c, p, thd):     @staticmethod class weight_quant(t.autograd.Function):     return (y - y_grad).detach() + y_grad     y_grad = x     y = x.round() def round_pass(x):      return (x - x_grad).detach() + x_grad, (y - y_grad).detach() + y_grad     y_grad = p * scale     x_grad = x * scale     scale = (1. - (p.detach() / c.detach() + 1e-12))     y = p     x = c def grad_p_scale(c, p):       return (y - y_grad).detach() + y_grad     y_grad = x * scale     y = x def grad_scale(x, scale):      return x def soft_pruner(x, block_size, p):  from .quantizer import Quantizer import math import torch as t ad  �              �  �  �  �  �  |  ^  <        �  �  �  �  m  %                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            plt.show()     plt.hist(module(x).flatten().detach()+0.1, bins = 400, alpha = 0.4)     module.hard_pruning = True     plt.hist(module(x).flatten().detach(), bins = 400)     plt.hist(x.flatten().detach(), bins = 400)          print(module(x))     print(x)          print(module.c, module.p)     module.p.data = t.tensor(0.4)     print(module.c, module.p)     module.init_from(x = x)     print(x)     x = t.randn((100,4,3,3))     module = SLsqQuan(bit = 8) if __name__ == "__main__": ''' ad     S     J       �  d  �  �  �  A  �  �  �  P    �  �  F  $  �  �  �  �  ^  A  �
  �
  `
  R
  
  �	  �	  �	  w	  L	  /	  �  �  M    	  �  �  J  �  �  >  �  �  c      �  �  �  �  �  ^  ]      �  �  �  �  R  ;  :  !  i  K  J  1  �  �  �  a  S  U                         else:             self.thd_pos = 2 ** bit - 1             self.thd_neg = 0             # unsigned activation is quantized to [0, 2^b-1]             assert not symmetric, "Positive quantization cannot be symmetric"         if all_positive:          super().__init__(bit)     def __init__(self, bit, all_positive=False, symmetric=True, per_channel=False, quant_mode = False, pruning_mode = False, block_size = 4, temperature = 1e-3, hard_pruning = False): class pqQuan(Quantizer):          return quant_x             #quant_x = (quant_x * mask - quant_x).detach() + quant_x             mask = self.soft_pruner(x, p_scale)         if (len(x.shape) == 4 and x.shape[1] != 1):          quant_x = quant_x * s          quant_x = (t.round(quant_x) - quant_x).detach() + quant_x          quant_x = t.clamp(quant_x, 0, self.thd_pos) * sign            quant_x = (x.abs() - p_scale) / s                  s = (c_scale - p_scale) / self.thd_pos         sign = x.sign()          #quant_x = self.weight_quantizer(x, c_scale, p_scale, self.thd_pos)         p_scale = grad_scale(self.p, p_grad_scale)         c_scale = grad_scale(self.c, c_grad_scale)             p_grad_scale = (self.thd_pos / x_numel) ** 0.5 * ((self.p+1e-20) / (self.c - self.p)).abs().detach() / 4             c_grad_scale = (self.thd_pos / x_numel) ** 0.5 / (self.c / (self.c - self.p)).detach() * self.thd_pos             x_numel = (x.abs() >= self.p).float().sum().detach()             #s_grad_scale = (x.abs().max().detach() / (self.thd_pos * x.numel())) ** 0.5             #s_grad_scale = 1.0 / ((x.numel()) ** 0.5)             #s_grad_scale = (self.thd_pos / x.numel()) ** 0.5 / 2             #s_grad_scale = 1.0 / ((self.thd_pos * x.numel()) ** 0.5)         else:             s_grad_scale = 1.0 / ((x.numel()) ** 0.5)             #s_grad_scale = (x.abs().max().detach() / (self.thd_pos * x.numel())) ** 0.5             #s_grad_scale = (self.thd_pos /  x.numel()) ** 0.5 / 2             #s_grad_scale = 1.0 / ((self.thd_pos * x.numel()) ** 0.5)         if self.per_channel:         self.p.data.clamp_(0.,self.c.data)     def forward(self, x):                  self.p = t.nn.Parameter(t.zeros([]))             self.c = t.nn.Parameter(s.clone().detach() * self.thd_pos)             s = x.detach().abs().mean() * 2 / (self.thd_pos ** 0.5)         else:             self.p = t.nn.Parameter(t.zeros_like(self.s))             self.c = t.nn.Parameter(s * self.thd_pos)             s = x.detach().abs().mean(dim = list(range(1, x.dim())), keepdim = True) * 2 / (self.thd_pos ** 0.5)         if self.per_channel:     def init_from(self, x, *args, **kwargs):          return hard_mask         hard_mask = hard_mask.repeat(1, self.block_size, 1, 1, 1).reshape(co,ci,kh,kw)         hard_mask = (score > 0).float()             return self.soft_mask             self.soft_mask = self.soft_mask.repeat(1, self.block_size, 1, 1, 1).reshape(co,ci,kh,kw)             self.soft_mask = _soft_mask             #_soft_mask = t.nn.functional.sigmoid(score)             _soft_mask = t.nn.functional.sigmoid(score/temperature)             #score = (score / temperature - score).detach() + score             #score = score - p             #p = grad_scale(p, p_grad_scale)             #p_grad_scale = temperature / ((self.c - self.p) * sigmoid_expectation).detach() / 2             #sigmoid_expectation = 1-t.nn.functional.sigmoid(-p / math.sqrt(1 + t.pi * temp_std ** 2 / 8)).detach()                          #temp_std = score.std().detach()             #temperature = (temp_score.abs().view(-1).sort()[0][int(score.numel()*self.temperature)] * 0.5).detach()             #temp_score = (score-p).detach()             temperature = (score.abs().view(-1).sort()[0][int(score.numel()*self.temperature)] * 0.5).detach() ad      �     c       �  �  �  z  [  Z  -    �  }  o      �  �  �  �  �  h  #    �  �  �  �  Q  7      
  �  \  >  5  
  �
  �
  �
  �
  b
  /
  
  �	  �	  �	  �	  	  ^	  ]	  <	  �  �  �  }  3    �  �  �  _    �  �  �  �  3  �  �  �  q  *  �  �  �  �  �  M  ?  �  �  �  z  `  W  ?    �  �  �  �  �  T  S  5  4    �  �  �              return quant_x             quant_x = quant_x * mask             mask = self.soft_pruner(x, p_scale)         if (len(x.shape) == 4):          quant_x = quant_x * s          quant_x = (t.round(quant_x) - quant_x).detach() + quant_x          quant_x = t.clamp(quant_x, 0, self.thd_pos) * sign            quant_x = (x.abs() - p_scale) / s                  s = (c_scale - p_scale + 1e-12) / self.thd_pos         sign = x.sign()                  #p_scale = self.p         #c_scale = self.c         p_scale = grad_scale(self.p, s_grad_scale)         c_scale = grad_scale(self.c, s_grad_scale)             s_grad_scale = 1.0 / ((self.thd_pos * x.numel()) ** 0.5)         else:             s_grad_scale = 1.0 / ((self.thd_pos * x.numel()) ** 0.5)         if self.per_channel:         self.p.data.clamp_(0.,self.c.data)     def forward(self, x):                  self.p = t.nn.Parameter(t.zeros([]))             self.c = t.nn.Parameter(s.clone().detach() * self.thd_pos)             s = x.detach().abs().mean() * 2 / (self.thd_pos ** 0.5)         else:             self.p = t.nn.Parameter(t.zeros_like(self.s))             self.c = t.nn.Parameter(s * self.thd_pos)             s = x.detach().abs().mean(dim = list(range(1, x.dim())), keepdim = True) * 2 / (self.thd_pos ** 0.5)         if self.per_channel:     def init_from(self, x, *args, **kwargs):          return hard_mask         hard_mask = hard_mask.repeat(1, self.block_size, 1, 1, 1).reshape(co,ci,kh,kw)         hard_mask = (score > 0).float()                      return _soft_mask             _soft_mask = _soft_mask.repeat(1, self.block_size, 1, 1, 1).reshape(co,ci,kh,kw)             self.soft_mask = _soft_mask             _soft_mask = t.nn.functional.sigmoid(score/ self.temperature)         if not self.hard_pruning:         score = x_reshape.abs().mean(dim = 1,keepdim = True).detach() - p          x_reshape = x.reshape(co // self.block_size, self.block_size, ci, kh, kw)         co, ci, kh, kw = x.shape      def soft_pruner(self, x, p):          self.temperature = temperature         self.hard_pruning = hard_pruning         self.mask_mean = 0.         self.block_size = block_size         self.soft_mask = None         self.weight_quantizer = weight_quant.apply         self.c = t.nn.Parameter(t.ones(1))         self.p= t.nn.Parameter(t.zeros(1))         self.per_channel = per_channel          self.thd_pos = 2 ** (bit - 1) - 1         self.thd_neg = -2 ** (bit - 1) + 1                  super().__init__(bit)     def __init__(self, bit, per_channel=False, symmetric = False, all_positive = False, hard_pruning = False, block_size = 4, temperature = 1e-3): class SLsqQuan(Quantizer): '''         return x         x = x * s_scale         x = round_pass(x)         x = t.clamp(x, self.thd_neg, self.thd_pos)         x = x / s_scale          s_scale = grad_scale(self.s, s_grad_scale)             s_grad_scale = 1.0 / ((self.thd_pos * x.numel()) ** 0.5)         else:             s_grad_scale = 1.0 / ((self.thd_pos * x.numel()) ** 0.5)         if self.per_channel:             self.init_mode = False             print(self.s)             self.init_from(x)         if self.init_mode:     def forward(self, x):              self.s = t.nn.Parameter(x.detach().abs().mean() * 2 / (self.thd_pos ** 0.5))         else:                 x.detach().abs().mean(dim=list(range(1, x.dim())), keepdim=True) * 2 / (self.thd_pos ** 0.5))             self.s = t.nn.Parameter(         if self.per_channel:     def init_from(self, x, *args, **kwargs):          self.init_mode = False         self.s = t.nn.Parameter(t.ones([]))         self.per_channel = per_channel                  self.thd_pos = 2 ** (bit - 1) - 1 ad  #   �     ]       �  �  _  -    �  �  h  g  @    �  �  �  �  z  \  7    �  �  �  �  w  	  �  �  h  .  -      �
  �
  �
  M
  
  �	  �	  �	  !	  �  �  �  w  ^  ]  C      �  �  �  d  H  )    �  �  �  t  <  *  �  �  �  p  o  O    �  �  �  �  �  �  O  1  0    �  �  o  G  '    �  �  x  F  4  �  �  �                                                     self.thd_neg = - 2 ** (bit - 1)                 # signed weight/activation is quantized to [-2^(b-1), 2^(b-1)-1]             else:                 self.thd_pos = 2 ** (bit - 1) - 1                 self.thd_neg = - 2 ** (bit - 1) + 1                 # signed weight/activation is quantized to [-2^(b-1)+1, 2^(b-1)-1]             if symmetric:         else:             print(self.thd_pos)             self.thd_pos = 2 ** bit - 1             self.thd_neg = 0             # unsigned activation is quantized to [0, 2^b-1]             assert not symmetric, "Positive quantization cannot be symmetric"         if all_positive:          super().__init__(bit)     def __init__(self, bit, all_positive=False, symmetric=True, per_channel=False): class LsqQuan(Quantizer):           return x_r             x_r = x_r * s_scale             x_r = round_pass(x_r)             x_r = t.clamp(x_r, self.thd_neg, self.thd_pos)             x_r = x_r / s_scale              s_scale = grad_scale(self.s, s_grad_scale)                  s_grad_scale = 1.0 / (x.numel() ** 0.5)                 #s_grad_scale = 1.0 / ((self.thd_pos * x.numel()) ** 0.5)             else:                 s_grad_scale = 1.0 / (x.numel() ** 0.5)                 #s_grad_scale = 1.0 / ((self.thd_pos * x.numel()) ** 0.5)             if self.per_channel:                  self.init_mode = False                 self.init_from(x)             if self.init_mode:         if self.quant_mode:                 x_r = x_r * mask                 mask = self.soft_pruner(x, self.p)             if (len(x.shape) == 4 and x.shape[1] != 1):         if self.pruning_mode:         x_r = x         self.p.data.clamp_(min = 0.)     def forward(self, x):          return hard_mask         hard_mask = hard_mask.repeat(1, self.block_size, 1, 1, 1).reshape(co,ci,kh,kw)         hard_mask = (score > 0).float()                      return self.soft_mask             self.soft_mask = self.soft_mask.repeat(1, self.block_size, 1, 1, 1).reshape(co,ci,kh,kw)             self.soft_mask = _soft_mask             _soft_mask = t.nn.functional.sigmoid(score/ self.temperature)         if not self.hard_pruning:         score = score / score.abs().max().detach()         score = x_reshape.abs().mean(dim = 1,keepdim = True).detach() - p          x_reshape = x.reshape(co // self.block_size, self.block_size, ci, kh, kw)         co, ci, kh, kw = x.shape      def soft_pruner(self, x, p):              self.p = t.nn.Parameter(t.zeros_like(self.s))             self.s = t.nn.Parameter(x.detach().abs().mean() * 2 / (self.thd_pos ** 0.5))         else:             self.s = t.nn.Parameter(t.zeros_like(self.s))                 x.detach().abs().mean(dim=list(range(1, x.dim())), keepdim=True) * 2 / (self.thd_pos ** 0.5))             self.s = t.nn.Parameter(         if self.per_channel:     def init_from(self, x, *args, **kwargs):          self.temperature = temperature         self.hard_pruning = hard_pruning         self.block_size = block_size         self.soft_mask = None         self.p= t.nn.Parameter(t.zeros([]))          self.pruning_mode = pruning_mode         self.quant_mode = quant_mode         self.init_mode = False         self.s = t.nn.Parameter(t.ones([]))         self.per_channel = per_channel                  self.thd_pos = 2 ** (bit - 1) - 1                 self.thd_neg = - 2 ** (bit - 1)                 # signed weight/activation is quantized to [-2^(b-1), 2^(b-1)-1]             else:                 self.thd_pos = 2 ** (bit - 1) - 1                 self.thd_neg = - 2 ** (bit - 1) + 1                 # signed weight/activation is quantized to [-2^(b-1)+1, 2^(b-1)-1]             if symmetric: 